newsp_inst : newsp PORT MAP (
		probe	 => probe_sig,
		source	 => source_sig
	);
