library verilog;
use verilog.vl_types.all;
entity sistema_completo_vlg_vec_tst is
end sistema_completo_vlg_vec_tst;
